/*
 *  This Verilog header file is where you can define or comment out areas
 *  during FPGA synthesis.
 */

`ifndef _ROBOCUP_HEADER_
`define _ROBOCUP_HEADER_

/**
 * Enable/Disable the module for the dribbler motor.
 */
`define DRIBBLER_MOTOR_EN


`endif  // _ROBOCUP_HEADER_
